<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-9.09313,14.8795,113.307,-45.6205</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>15.5,-12.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>13.5,-8</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>14,-18</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>59.5,-9.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>60,-16</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>BA_NAND2</type>
<position>28.5,-8.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>28.5,-17</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>BA_NAND2</type>
<position>40.5,-9.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND2</type>
<position>40.5,-16</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-16,24,-9.5</points>
<intersection>-16 3</intersection>
<intersection>-12.5 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-9.5,25.5,-9.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-12.5,24,-12.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-16,25.5,-16</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-8,25.5,-8</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>25.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>25.5,-8,25.5,-7.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-8 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-12,58.5,-12</points>
<intersection>35.5 6</intersection>
<intersection>43.5 7</intersection>
<intersection>58.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>35.5,-15,35.5,-12</points>
<intersection>-15 9</intersection>
<intersection>-12 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>43.5,-12,43.5,-9.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>-12 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>58.5,-12,58.5,-9.5</points>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>35.5,-15,37.5,-15</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>35.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-13.5,59,-13.5</points>
<intersection>37.5 3</intersection>
<intersection>43.5 5</intersection>
<intersection>59 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-13.5,37.5,-10.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>59,-16,59,-13.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>43.5,-16,43.5,-13.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-17,37.5,-17</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-8.5,37.5,-8.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-18,25.5,-18</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 9></circuit>